../calculator/bcd_mux.sv