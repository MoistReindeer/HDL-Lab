../calculator/display.sv