../calculator/seg_dec.sv